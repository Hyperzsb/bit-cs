module pow3 (
    input[2:0] in,
    output[5:0] out
);

assign out = in * in;

endmodule // 